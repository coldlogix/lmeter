LPIC3 9 32 0.197000
LCP2 27 13 0.031000
LPJC2 0 10 0.034000
LPJC3 29 0 0.027000
LPJC1 38 0 0.024000
LPIC1 21 36 0.327000
LPDA 33 17 0.371000
LPJDA1 0 18 0.035000
LPJDA2 0 14 0.015000
LPJA1 12 0 0.018000
LPIA1 25 39 0.248000
LPJA2 0 34 0.021000
LPIA2 35 28 0.744000
LPJA4 0 31 0.045000
LPIA3 4 1 0.216000
LPIC2 27 30 0.544000
LPIDA 23 22 0.345000
LPJA3 26 0 0.030000
LDAQ 23 33 2.067000
IC3 9 0 1.330000
IC1 36 0 3.210000
IDA 22 0 0.770000
IA3 1 0 2.190000
IA2 28 0 1.030000
IC2 30 0 2.650000
IA1 39 0 1.100000
LC2 7 13 0.467000
LC4 32 20 0.104000
LC3 7 32 0.294000
LC1 7 21 0.329000
LCIN 2 21 0.111000
LXA2 4 5 0.752000
LXA1 4 19 0.391000
LA4 19 37 0.673000
L6 8 27 0.120000
LA2 16 25 0.376000
LAOUT 3 35 0.489000
LA5 19 35 0.603000
LA1 33 16 0.422000
LAIN 6 23 0.277000
LCOUT 11 8 0.528000
LA3 25 37 0.754000
LCDA 17 15 0.488000
JC3 32 29 2.680000
JC2 13 10 2.930000
JC1 21 38 3.460000
JA4 4 31 1.780000
JA2 37 34 2.210000
JA1 16 12 2.440000
JA3 35 26 1.780000
JDA2 17 14 1.580000
JDA1 23 18 2.680000
JDA3 8 15 2.440000
PCLKOUT 11 0 1.0
PAOUT 3 0 1.0
PAIN 6 0 1.0
PCLKOUT2 20 0 1.0
PAOUT2 5 0 1.0
PCLKIN 2 0 1.0
.END
