KX LJ6 LJ1 0.0
K1 L17 L10 0.0860
K2 L7 L8 0.0490
K3 L26 L17 0.0170
K4 L3 L1 0.0140
L11 12 11 0.046000
L22 19 9 0.082000
LJ2 8 0 0.049000
LJ1 5 0 0.037000
LJ3 21 0 0.059000
LJ6 22 0 0.045000
L10 13 6 0.570000
L25 19 7 0.149000
L12 23 7 0.307000
L9 16 10 0.248000
J13 9 0 1.490000
J1 3 5 2.010000
J2 2 8 2.010000
J3 18 21 2.010000
J4 12 22 2.600000
L17 7 14 0.819000
L4 2 18 1.511000
L2 3 10 0.746000
L3 10 2 0.754000
L1 3 1 0.550000
L5 6 18 0.781000
L6 11 6 0.532000
L7 4 12 0.889000
L8 20 11 0.657000
L26 17 19 1.593000
I3 23 0 1.190000
IC1 16 0 2.800000
IC2 13 0 3.100000
RJ2 0 2 0.300000
RJ3 0 18 0.300000
RJ6 0 12 0.300000
PSI 14 0 1.0
PSO 17 0 1.0
PCLMO 20 0 1.0
PCLMI 1 0 1.0
PNRO 4 0 1.0
.END
